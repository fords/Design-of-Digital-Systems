//Verilog HDL for "zxw_lib", "zxw_inv3" "test"


module zxw_inv3 ( );

endmodule
