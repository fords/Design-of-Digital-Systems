//Verilog HDL for "zxw_lib", "zxw_inv4" "zxw_inv4Verilog"


module zxw_inv4 (in1,out1
);

	input in1;
	output out1;
	not (out1,in1);
endmodule
