*
*
*
*                       LINUX           Fri Oct 31 22:57:03 2014
*
*
*
*  PROGRAM  advgen
*
*  CDL LIBRARY
*
*
*

*
.SUBCKT zxw_dff gnd! D Q Qbar phi1 phi2
*
*
*  caps2d version: 7
*
*
*       TRANSISTOR CARDS
*
*
M50	net0183#2	net0346#4	net0268	gnd!#1	nmos	L=0.6
+ W=4.8
+ AD=6.57	AS=3.765	PD=8	PS=1.8
M51	net0268	net076#4	gnd!#16	gnd!#1	nmos	L=0.6
+ W=4.8
+ AD=3.765	AS=3.765	PD=1.8	PS=1.8
M49	net0260	phi1#5	gnd!#16	gnd!#1	nmos	L=0.6	W=4.8
+ AD=3.765	AS=3.765	PD=1.8	PS=1.8
M48	net0183#3	net0130#6	net0260	gnd!#1	nmos	L=0.6
+ W=4.8
+ AD=6.57	AS=3.765	PD=8	PS=1.8
M10	net076#7	phi1#4	gnd!#15	gnd!#1	nmos	L=0.6	W=2.4
+ AD=4	AS=2.24	PD=6.6	PS=2.3
M36	net0255#2	net0183#11	gnd!#15	gnd!#1	nmos	L=0.6
+ W=2.4
+ AD=4	AS=2.24	PD=6.6	PS=2.3
M27	net0261#3	net0255#8	gnd!#14	gnd!#1	nmos	L=0.6
+ W=2.4
+ AD=4.11	AS=2.295	PD=6.8	PS=2.4
M26	net0346#7	net0261#8	gnd!#14	gnd!#1	nmos	L=0.6
+ W=2.4
+ AD=4.11	AS=2.295	PD=6.8	PS=2.4
M31	Q#3	net0261#11	gnd!#13	gnd!#1	nmos	L=0.6	W=2.4
+ AD=4.11	AS=2.295	PD=6.8	PS=2.4
M30	Qbar#3	net0255#6	gnd!#13	gnd!#1	nmos	L=0.6	W=2.4
+ AD=4.11	AS=2.295	PD=6.8	PS=2.4
M45	net0187#2	net0286#4	net0216	gnd!#1	nmos	L=0.6
+ W=4.8
+ AD=6.57	AS=3.765	PD=8	PS=1.8
M46	net0216	net0220#4	gnd!#12	gnd!#1	nmos	L=0.6
+ W=4.8
+ AD=3.765	AS=3.765	PD=1.8	PS=1.8
M44	net0208	phi2#6	gnd!#12	gnd!#1	nmos	L=0.6	W=4.8
+ AD=3.765	AS=3.765	PD=1.8	PS=1.8
M43	net0187#3	net0211#3	net0208	gnd!#1	nmos	L=0.6
+ W=4.8
+ AD=6.57	AS=3.765	PD=8	PS=1.8
M20	net0211#6	D#4	gnd!#19	gnd!#1	nmos	L=0.6	W=2.4
+ AD=4	AS=4	PD=6.6	PS=6.6
M47	net0220#7	phi2#4	gnd!#18	gnd!#1	nmos	L=0.6	W=2.4
+ AD=4	AS=2.24	PD=6.6	PS=2.3
M34	net0132	net0187#10	gnd!#18	gnd!#1	nmos	L=0.6
+ W=2.4
+ AD=4	AS=2.24	PD=6.6	PS=2.3
M22	net0130#3	net0132#6	gnd!#17	gnd!#1	nmos	L=0.6
+ W=2.4
+ AD=4.11	AS=2.295	PD=6.8	PS=2.4
M24	net0286#7	net0130#10	gnd!#17	gnd!#1	nmos	L=0.6
+ W=2.4
+ AD=4.11	AS=2.295	PD=6.8	PS=2.4
M53	net0339	net0346#3	vdd!#16	vdd!#2	pmos	L=0.6
+ W=9.6
+ AD=12.48	AS=7.2	PD=12.2	PS=1.5
M54	net0339#3	net076#3	vdd!#16	vdd!#2	pmos	L=0.6
+ W=9.6
+ AD=7.2	AS=7.2	PD=1.5	PS=1.5
M55	net0183#7	phi1#7	net0339#3	vdd!#2	pmos	L=0.6	W=9.6
+ AD=7.2	AS=7.2	PD=1.5	PS=1.5
M52	net0183#7	net0130#7	net0339#5	vdd!#2	pmos	L=0.6
+ W=9.6
+ AD=7.2	AS=12.48	PD=1.5	PS=12.2
M15	net076#5	phi1#6	vdd!#15	vdd!#2	pmos	L=0.6	W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M37	net0255	net0183#8	vdd!#15	vdd!#2	pmos	L=0.6
+ W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M29	net0261	net0255#9	vdd!#14	vdd!#2	pmos	L=0.6
+ W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M28	net0346#5	net0261#6	vdd!#14	vdd!#2	pmos	L=0.6
+ W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M32	Q#4	net0261#9	vdd!	vdd!#2	pmos	L=0.6	W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M33	Qbar#1	net0255#5	vdd!	vdd!#2	pmos	L=0.6	W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M39	net0283	net0286#3	vdd!#13	vdd!#2	pmos	L=0.6
+ W=9.6
+ AD=12.48	AS=7.2	PD=12.2	PS=1.5
M40	net0283#3	net0220#3	vdd!#13	vdd!#2	pmos	L=0.6
+ W=9.6
+ AD=7.2	AS=7.2	PD=1.5	PS=1.5
M41	net0187#7	phi2#7	net0283#3	vdd!#2	pmos	L=0.6	W=9.6
+ AD=7.2	AS=7.2	PD=1.5	PS=1.5
M38	net0187#7	net0211#4	net0283#5	vdd!#2	pmos	L=0.6
+ W=9.6
+ AD=7.2	AS=12.48	PD=1.5	PS=12.2
M21	net0211#5	D#5	vdd!#19	vdd!#2	pmos	L=0.6	W=4.8
+ AD=6.79	AS=6.9	PD=8.4	PS=8.6
M42	net0220#6	phi2#3	vdd!#18	vdd!#2	pmos	L=0.6	W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M35	net0132#3	net0187#12	vdd!#18	vdd!#2	pmos	L=0.6
+ W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M23	net0130	net0132#5	vdd!#17	vdd!#2	pmos	L=0.6
+ W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
M25	net0286#5	net0130#8	vdd!#17	vdd!#2	pmos	L=0.6
+ W=4.8
+ AD=6.79	AS=3.875	PD=8.4	PS=2
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Re1	net0286#3	net0286#2	  337.2261
Re2	net0286#2	net0286#4	  211.6161
Re3	net0220#3	net0220#2	  360.5432
Re4	net0220#2	net0220#4	  171.6105
Re5	net0211	net0211#2	  340.8918
Re6	net0211#2	net0211#3	  213.1135
Re7	net0211#2	net0211#4	  385.2272
Re8	D#1	D#4	  232.2549
Re9	D#4	D#5	  600.5174
Re10	phi2#3	phi2#4	  596.9937
Re11	phi2#4	phi2#5	  125.2420
Re12	phi2#5	phi2#6	  871.5280
Re13	phi2#5	phi2#2	   13.5000
Re14	phi2#6	phi2#7	  570.8168
Re15	net0187#10	net0187#11	  405.8915
Re16	net0187#11	net0187#8	   10.5000
Re17	net0187#11	net0187#12	  196.3821
Re18	net0132#5	net0132#6	  605.0000
Re19	net0132#6	net0132#4	  226.3773
Re20	net0346#3	net0346#2	  335.5503
Re21	net0346#2	net0346#4	  209.3938
Re22	net076#3	net076#2	  361.2143
Re23	net076#2	net076#4	  171.2626
Re24	net0130#6	net0130#7	  598.5237
Re25	net0130#7	net0130#8	 1070.2894
Re26	net0130#8	net0130#9	  186.6294
Re27	net0130#9	net0130#5	   11.0526
Re28	net0130#9	net0130#10	  414.1294
Re29	phi1#2	phi1#3	   15.0000
Re30	phi1#3	phi1#4	  122.5443
Re31	phi1#4	phi1#5	  771.5276
Re32	phi1#3	phi1#6	  472.5443
Re33	phi1#5	phi1#7	  570.8168
Re34	net0183#8	net0183#9	  195.2420
Re35	net0183#9	net0183#10	   49.0000
Re36	net0183#9	net0183#11	  405.2420
Re37	net0261#6	net0261#7	  478.0177
Re38	net0261#7	net0261#5	   11.6667
Re39	net0261#7	net0261#8	  123.0177
Re40	net0261#9	net0261#10	  467.5000
Re41	net0261#10	net0261#11	  112.5000
Re42	net0255#5	net0255#6	  605.0000
Re43	net0255#6	net0255#7	  408.3697
Re44	net0255#7	net0255#4	  101.0413
Re45	net0255#7	net0255#8	  124.2649
Re46	net0255#8	net0255#9	  605.0000
Rc1	net0187	net0187#2	   17.1889
Rc2	net0286	net0286#2	   41.0000
Rc3	net0283	net0283#2	   12.3944
Rc4	net0220	net0220#2	   41.0000
Rc5	net0283#3	net0283#4	   12.3944
Rc6	net0187#4	net0187#5	    0.8760
Rc7	net0187#4	net0187#6	    1.1889
Rc8	net0187#5	net0187#7	   11.3000
Rc9	net0187#3	net0187#4	   16.0000
Rc10	net0283#5	net0283#6	   12.3944
Rc11	net0211#5	net0211#7	   21.1816
Rc12	net0211#7	net0211	    0.2419
Rc13	net0211#6	net0211#7	   26.6667
Rc14	D#1	D#2	   20.5000
Rc15	net0220#5	net0220#6	   20.8932
Rc16	net0220#5	net0220#7	   26.9169
Rc17	phi2#1	phi2#2	   41.0000
Rc18	net0187#8	net0187#9	   41.0000
Rc19	net0132#2	net0132#3	   21.1435
Rc20	net0132#2	net0132#4	   40.2597
Rc21	net0132	net0132#2	   26.6667
Rc22	net0130	net0130#2	   20.3589
Rc23	net0130#2	net0130#3	   27.4506
Rc24	net0130#4	net0130#5	   41.0000
Rc25	net0286#5	net0286#6	   20.7272
Rc26	net0286#6	net0286#7	   27.0822
Rc27	net0183	net0183#2	   17.1889
Rc28	net0346	net0346#2	   41.0000
Rc29	net0339	net0339#2	   12.3944
Rc30	net076	net076#2	   41.0000
Rc31	net0339#3	net0339#4	   12.3944
Rc32	net0183#4	net0183#5	    0.8760
Rc33	net0183#4	net0183#6	    1.1889
Rc34	net0183#5	net0183#7	   11.3000
Rc35	net0183#3	net0183#4	   16.0000
Rc36	net0339#5	net0339#6	   12.3944
Rc37	net076#5	net076#6	   20.8925
Rc38	net076#6	net076#7	   26.9169
Rc39	phi1#1	phi1#2	   41.0000
Rc40	net0183#10	net0183#12	    1.0000
Rc41	net0255	net0255#3	   21.1428
Rc42	net0255#3	net0255#4	   40.2597
Rc43	net0255#2	net0255#3	   26.6667
Rc44	net0261	net0261#2	   20.9067
Rc45	net0261#2	net0261#3	   26.9028
Rc46	net0261#4	net0261#5	   41.0000
Rc47	net0346#5	net0346#6	   20.7367
Rc48	net0346#6	net0346#7	   27.0728
Rc49	Q#1	Q#2	    0.5216
Rc50	Q#2	Q#3	   27.2761
Rc51	Q#2	Q#4	   20.4347
Rc52	net0261#12	net0261#10	   41.0000
Rc53	Qbar#1	Qbar#2	   20.4316
Rc54	Qbar#2	Qbar#3	   27.2930
Rc55	gnd!#1	gnd!#2	    5.9194
Rc56	gnd!#2	gnd!#3	9.040E-02
Rc57	gnd!#3	gnd!#4	8.757E-02
Rc58	gnd!#4	gnd!#5	1.970E-02
Rc59	gnd!#5	gnd!#6	    0.1196
Rc60	gnd!#6	gnd!#7	    0.1150
Rc61	gnd!#7	gnd!#8	1.085E-02
Rc62	gnd!#8	gnd!#9	8.757E-02
Rc63	gnd!#9	gnd!#10	8.119E-02
Rc64	gnd!#10	gnd!#11	6.185E-02
Rc65	gnd!#11	gnd!	1.947E-02
Rc66	gnd!	gnd!#12	   16.3788
Rc67	gnd!#2	gnd!#13	   27.1041
Rc68	gnd!#3	gnd!#14	   27.1041
Rc69	gnd!#4	gnd!#15	   27.0994
Rc70	gnd!#6	gnd!#16	   16.3477
Rc71	gnd!#8	gnd!#17	   27.1041
Rc72	gnd!#9	gnd!#18	   27.0994
Rc73	gnd!#10	gnd!#19	   27.0994
Rc74	gnd!#1	gnd!#5	    6.2500
Rc75	gnd!#1	gnd!#7	    5.8824
Rc76	gnd!#1	gnd!#11	    5.8824
Rc77	vdd!	vdd!#3	   20.3656
Rc78	vdd!#3	vdd!#4	6.787E-02
Rc79	vdd!#4	vdd!#5	8.757E-02
Rc80	vdd!#5	vdd!#6	6.362E-02
Rc81	vdd!#6	vdd!#7	8.416E-02
Rc82	vdd!#7	vdd!#8	    0.1173
Rc83	vdd!#8	vdd!#9	1.758E-02
Rc84	vdd!#9	vdd!#10	7.070E-02
Rc85	vdd!#10	vdd!#11	7.269E-02
Rc86	vdd!#11	vdd!#12	7.637E-02
Rc87	vdd!#12	vdd!#13	   11.7095
Rc88	vdd!#4	vdd!#14	   20.3524
Rc89	vdd!#5	vdd!#15	   20.3571
Rc90	vdd!#7	vdd!#16	   11.6571
Rc91	vdd!#8	vdd!#17	   20.3524
Rc92	vdd!#10	vdd!#18	   20.3571
Rc93	vdd!#11	vdd!#19	   20.3571
Rc94	vdd!#2	vdd!#3	    5.3333
Rc95	vdd!#2	vdd!#6	    5.0000
Rc96	vdd!#2	vdd!#9	    5.3333
Rc97	vdd!#2	vdd!#12	    5.0000
Rb1	net0187#6	net0187	    0.7933
Rb2	net0283#6	net0283#4	    0.3967
Rb3	net0283#4	net0283#2	    0.3967
Rb4	D#2	D	    0.5000
Rb5	net0220#5	net0220	    2.2750
Rb6	phi2#1	phi2	    1.0000
Rb7	net0187#9	net0187#5	    2.1144
Rb8	net0130#4	net0130#2	    1.2361
Rb9	net0286#6	net0286	    3.5358
Rb10	net0183#6	net0183	    0.7933
Rb11	net0339#6	net0339#4	    0.3967
Rb12	net0339#4	net0339#2	    0.3967
Rb13	net076#6	net076	    1.7886
Rb14	phi1#1	phi1#8	    1.0000
Rb15	net0183#12	net0183#5	    1.6328
Rb16	net0346#6	net0346	    3.0447
Rb17	Q#1	Q	    0.5000
Rb18	net0261#12	net0261#4	    0.5100
Rb19	net0261#4	net0261#2	    1.2361
Rb20	Qbar#2	Qbar	    1.0000
Ra3	phi1	phi1#8	3.250E-02
*
*       CAPACITOR CARDS
*
*
C1	net0183#6	gnd!#16	7.650E-17
C2	vdd!#19	D#5	1.631E-16
C3	net0187#5	vdd!#19	1.374E-17
C4	vdd!#7	net0130#7	2.061E-16
C5	vdd!#19	net0220#6	7.913E-17
C6	net0339#4	net0183#7	7.312E-17
C7	net076#5	net0130#7	1.159E-17
C8	net0183#7	net0339#5	1.758E-16
C9	net0346#5	vdd!#2	3.141E-17
C10	net0187#6	phi2#6	2.350E-17
C11	vdd!#17	net0130#5	1.454E-17
C12	Q#3	Qbar#3	6.721E-18
C13	gnd!#12	net0286#4	8.334E-17
C14	Q#1	net0261#9	1.456E-16
C15	net0130#3	net0132#6	2.037E-16
C16	net0211#5	D#5	2.733E-16
C17	gnd!#8	net0130#10	2.476E-17
C18	net0130#10	gnd!#1	5.688E-16
C19	net0339#3	net0183#5	1.527E-16
C20	net0187#5	net0211#4	9.616E-17
C21	phi2#6	net0211#2	2.380E-17
C22	phi1#3	gnd!#1	4.207E-16
C23	gnd!#14	net0261#4	9.608E-17
C24	Q	net0261#9	1.037E-17
C25	net0339#5	net0130#7	2.701E-16
C26	D	net0211#4	1.075E-16
C27	net0255#2	net0183#11	1.827E-16
C28	Q	net0261#6	9.814E-18
C29	Q#1	Qbar#2	1.697E-16
C30	vdd!#2	net0132#5	7.193E-17
C31	net0187#5	net0211#5	1.165E-16
C32	net0283#5	D#5	1.107E-17
C33	net076#2	phi1#7	3.298E-17
C34	net0346#6	phi1#3	4.239E-17
C35	Q	net0255#6	3.441E-17
C36	phi1	net0255#9	1.830E-17
C37	net0183#7	net0130#7	1.580E-16
C38	net0187#5	phi2#7	1.492E-16
C39	net0261#12	Q#1	2.165E-17
C40	net0132#6	gnd!#1	6.147E-16
C41	net0211#5	net0220#6	1.027E-17
C42	gnd!#15	net0183#11	9.678E-17
C43	phi2#2	gnd!#1	2.078E-16
C44	net0130#3	net0187#10	9.317E-18
C45	phi1#8	net0255#2	5.728E-17
C46	Q	net0261#10	3.137E-17
C47	D	net0286#6	1.143E-16
C48	net076#6	net0130#6	2.324E-17
C49	D	net0187#9	1.288E-16
C50	D	phi2#1	2.055E-17
C51	net0283#4	phi2#7	2.079E-17
C52	D	net0220#5	1.448E-16
C53	net0283#6	net0187#7	7.887E-17
C54	net0339#3	net0130#7	1.123E-17
C55	net0283#3	net0187#7	1.758E-16
C56	gnd!#6	net0183#6	1.909E-16
C57	net0346#6	net0183#9	3.695E-17
C58	vdd!#7	phi1#7	1.421E-17
C59	net0339#5	phi1#7	4.846E-18
C60	net0255#2	net0261#3	1.452E-16
C61	net0187#5	net0211#6	2.929E-17
C62	net0283#3	net0220#2	3.940E-17
C63	D	gnd!#1	8.810E-17
C64	net0346#7	net0255#7	3.239E-17
C65	Q	Qbar#2	4.157E-17
C66	Q	net0261#12	1.204E-16
C67	Q	net0346#6	3.878E-17
C68	gnd!#17	net0132#4	3.319E-17
C69	net0132#5	net0130#9	3.999E-17
C70	net0255#7	net0261#8	4.980E-17
C71	net0286#5	vdd!#8	1.213E-16
C72	net0339#4	vdd!#2	2.941E-17
C73	net0346#6	net0255#2	1.306E-16
C74	Q#3	gnd!#13	9.829E-17
C75	net0132#3	net0130#2	1.813E-16
C76	net0183#7	phi1#7	1.513E-16
C77	net0220#7	phi2#5	2.509E-17
C78	net0283#5	net0211#4	2.443E-16
C79	net0187#10	gnd!#1	4.902E-16
C80	net0183#6	net0130#6	5.664E-17
C81	gnd!#12	net0220#2	4.927E-17
C82	D#1	gnd!#1	8.029E-16
C83	phi1#4	net0183#11	1.163E-17
C84	net0283#4	net0220#3	2.306E-17
C85	gnd!#15	phi1#4	1.042E-16
C86	D	net0220#7	2.216E-17
C87	D	net0220#6	7.425E-17
C88	D	gnd!#19	4.368E-17
C89	D	vdd!#19	7.618E-17
C90	D	net0211#5	3.684E-17
C91	D	net0211#6	1.730E-17
C92	net0187#5	net0283#5	2.348E-16
C93	Q#1	net0346#6	2.216E-17
C94	net0339#3	phi1#7	2.773E-16
C95	net0255#8	net0261#7	4.864E-17
C96	net0187#5	net0283#6	3.441E-17
C97	net0183#5	net0130#6	1.210E-17
C98	D	net0211#2	3.183E-17
C99	Q	gnd!#1	7.546E-17
C100	Q	Qbar#1	1.884E-17
C101	gnd!#14	net0261#7	1.765E-17
C102	Q	vdd!#2	2.889E-16
C103	Q	Qbar#3	1.779E-17
C104	gnd!#18	net0187#10	9.682E-17
C105	net0283#5	vdd!#2	1.144E-16
C106	Q	gnd!#13	7.607E-17
C107	net0187#7	net0211#4	1.520E-16
C108	net0286#7	gnd!#1	5.492E-17
C109	gnd!#15	net0255#4	4.048E-17
C110	Q	net0346#5	5.487E-18
C111	net0346#6	net0261#7	1.972E-16
C112	net0339#4	vdd!#16	8.058E-17
C113	vdd!#13	net0220#2	8.773E-17
C114	Q	vdd!#14	5.546E-18
C115	Q	gnd!#14	1.245E-17
C116	phi1#3	net0183#11	5.365E-17
C117	net0183#6	phi1#5	2.351E-17
C118	net0130#3	net0132#4	3.206E-17
C119	D	gnd!#10	3.676E-16
C120	net0286#6	net0346#2	2.593E-17
C121	phi2#4	gnd!#1	4.049E-16
C122	net0261#7	gnd!#1	2.578E-16
C123	phi1	net0346#6	1.504E-16
C124	D	vdd!#11	3.522E-16
C125	net076#7	phi1#4	1.458E-16
C126	vdd!#7	net076#3	5.994E-17
C127	phi1#8	gnd!#15	9.603E-17
C128	phi1#8	gnd!#4	5.161E-16
C129	phi1	net0183#12	1.378E-16
C130	net076#7	gnd!#4	1.427E-17
C131	net0187#9	net0132#3	2.032E-17
C132	phi1	net076#6	2.880E-17
C133	net0183#10	vdd!#15	4.928E-17
C134	net0283#3	net0211#4	4.538E-18
C135	net0283#5	phi2#7	5.034E-18
C136	net0346#6	Q#2	1.692E-16
C137	net0220#2	phi2#6	7.609E-17
C138	net0132#5	net0130#5	3.141E-17
C139	net0183#12	phi1#6	3.022E-17
C140	net0339#3	net076#3	2.121E-16
C141	gnd!#3	net0346#7	3.549E-17
C142	net0261#4	net0346#6	2.412E-16
C143	net0211#6	gnd!#19	1.043E-16
C144	net0211#5	vdd!#19	1.866E-16
C145	net0286#6	net0130#9	1.602E-16
C146	gnd!#9	net0187#10	2.533E-17
C147	net0283#2	net0286#3	2.306E-17
C148	phi1#5	net0130#6	7.383E-17
C149	gnd!#18	phi2#4	7.871E-17
C150	D#4	gnd!#1	4.444E-16
C151	net0346#5	Q#4	1.664E-16
C152	net0187#7	phi2#7	1.513E-16
C153	net0255#2	net0261#2	1.647E-16
C154	net0220#2	gnd!#1	4.182E-16
C155	gnd!#9	phi2#1	9.768E-17
C156	vdd!#13	net0286#2	5.016E-17
C157	Q	net0261#7	1.887E-17
C158	vdd!#16	net076#3	2.148E-16
C159	Q	gnd!#2	3.273E-16
C160	phi2#5	D#1	1.832E-17
C161	gnd!#9	phi2#5	2.746E-16
C162	phi1#8	gnd!#1	7.363E-17
C163	net0346#6	net0261#2	2.370E-16
C164	net076#5	net0183#10	2.140E-17
C165	net0339#3	net0183#7	1.758E-16
C166	vdd!#2	net0211#4	5.207E-17
C167	net0255#2	gnd!#1	8.802E-17
C168	net0346#2	net076#2	8.395E-17
C169	net0187#7	vdd!#2	1.144E-16
C170	gnd!#18	net0132#4	4.220E-17
C171	net076#4	phi1#5	1.789E-17
C172	gnd!#14	net0255#7	8.086E-17
C173	net0283#3	phi2#7	2.773E-16
C174	net0187#8	net0132#3	2.221E-16
C175	vdd!#7	net0346#3	6.035E-17
C176	net0339#3	net0346#3	4.497E-18
C177	net0220#7	phi2#4	8.294E-17
C178	net0211#3	gnd!#1	3.858E-16
C179	net0255#7	gnd!#1	1.110E-15
C180	phi1#8	net076#7	1.047E-16
C181	net0183#3	net0130#6	3.161E-16
C182	net0286#2	gnd!#1	3.527E-16
C183	net0339#6	net0130#7	1.606E-17
C184	net0346#6	net0183#12	9.615E-17
C185	phi1	net0255#2	1.611E-17
C186	net0261#9	net0255#5	3.948E-17
C187	Q#2	net0261#9	5.657E-17
C188	net0339#2	vdd!#16	9.422E-17
C189	net0187#5	net0283#4	1.162E-17
C190	phi1	vdd!#15	1.035E-16
C191	net0286#6	gnd!#1	2.648E-17
C192	phi1	net076#5	8.540E-17
C193	vdd!#18	net0132#3	1.849E-16
C194	net0187#6	gnd!#12	1.393E-16
C195	net0286#6	net0187#8	4.708E-17
C196	phi2#3	net0187#8	9.601E-17
C197	vdd!#16	net0346#3	2.069E-16
C198	net0283#4	net0187#7	7.252E-17
C199	vdd!#2	phi2#7	4.946E-17
C200	Q#2	Qbar#1	5.929E-18
C201	net0346#4	net076#4	2.204E-17
C202	net0183#5	net0130#7	1.512E-16
C203	net0220#6	vdd!#10	9.295E-17
C204	net0255#6	net0261#10	6.561E-17
C205	net0187#9	vdd!#18	4.600E-17
C206	phi1#1	net0346#6	9.413E-17
C207	vdd!#13	gnd!#1	6.208E-17
C208	gnd!#10	phi2#5	3.604E-16
C209	gnd!#15	net0255#2	1.246E-16
C210	net0283#3	net0187#5	1.576E-16
C211	net0183#12	vdd!#15	3.519E-17
C212	phi2#6	gnd!#1	1.581E-15
C213	net0255#9	net0261#6	5.105E-17
C214	net0346#7	Q#3	1.419E-16
C215	gnd!#4	net0183#11	2.257E-17
C216	net0283#3	net0220#3	2.121E-16
C217	phi2#1	gnd!#18	4.947E-17
C218	phi1#5	net0183#3	8.114E-17
C219	phi1#1	net0255#2	4.592E-17
C220	vdd!#17	net0286#5	1.849E-16
C221	net0183#5	phi1#7	1.476E-16
C222	vdd!#7	net0130#8	2.881E-16
C223	net0346#6	net076#6	1.348E-16
C224	Qbar#2	net0261#10	9.848E-18
C225	net0255#2	net0183#9	6.096E-17
C226	net0187#8	vdd!#18	8.261E-17
C227	net0130#3	gnd!#1	6.802E-17
C228	net0339#4	phi1#7	2.305E-17
C229	net0283#3	vdd!#2	5.088E-17
C230	vdd!#8	net0130#8	3.502E-16
C231	Qbar#1	net0255#5	1.834E-16
C232	vdd!#13	net0220#3	2.777E-16
C233	net0220#4	gnd!#1	3.588E-16
C234	phi1#8	net0346#6	2.122E-17
C235	phi1#8	net0183#3	2.704E-17
C236	vdd!#13	net0283#3	3.683E-16
C237	phi1#6	net0183#8	1.736E-17
C238	net0261#12	gnd!#1	7.830E-17
C239	gnd!#19	D#4	1.114E-16
C240	net0183#12	net076#5	1.206E-16
C241	net0286#6	net0130#4	4.843E-17
C242	net076#6	net0255#2	1.269E-17
C243	net0132#6	net0130#10	4.659E-17
C244	net0339#4	net076#3	2.306E-17
C245	net0187#9	net0220#6	1.177E-16
C246	net0339#3	phi1#5	5.674E-18
C247	Q#1	net0261#10	1.312E-16
C248	net0283#3	net0286#3	4.497E-18
C249	gnd!#4	phi1#4	1.873E-16
C250	net0255#6	gnd!#1	1.280E-15
C251	phi1#1	gnd!#15	9.225E-17
C252	net0255#8	net0261#5	2.585E-17
C253	Qbar#1	net0261#9	6.220E-18
C254	net0283#5	net0211#5	3.250E-16
C255	net0220#6	net0187#8	3.137E-17
C256	net0261#3	net0255#7	4.005E-17
C257	net0286#5	net0130#8	1.418E-16
C258	net0286#4	gnd!#1	4.393E-16
C259	net0339#3	vdd!#7	1.144E-16
C260	net0220#6	net0132#3	1.376E-17
C261	phi2#1	net0220#7	8.201E-17
C262	gnd!#16	phi1#5	1.454E-16
C263	phi1	vdd!#5	4.951E-16
C264	vdd!#2	net0261#9	5.470E-17
C265	net0255#9	net0261#7	2.373E-17
C266	phi1#7	net0130#7	4.516E-17
C267	vdd!#15	net0183#9	3.205E-17
C268	net076#5	vdd!#15	1.600E-16
C269	net0283#5	net0211#2	2.646E-17
C270	net0286#6	net0130#2	1.029E-16
C271	vdd!#14	net0346#5	1.849E-16
C272	D#2	gnd!#10	3.278E-17
C273	gnd!#9	net0220#7	1.695E-17
C274	vdd!#13	net0286#3	2.700E-16
C275	net076#6	phi1#3	1.604E-16
C276	net076#3	net0130#7	2.568E-17
C277	net0286#6	net0130#10	4.552E-17
C278	vdd!#17	net0130#8	1.196E-16
C279	net076#7	gnd!#1	2.070E-16
C280	vdd!#8	net0132#5	1.298E-17
C281	net0220#5	net0187#8	7.818E-18
C282	gnd!#15	phi1#3	3.026E-17
C283	phi2#2	net0220#7	1.972E-17
C284	net076#3	phi1#7	1.826E-17
C285	net0220#2	phi2#7	3.220E-17
C286	net0211#6	D#4	2.847E-16
C287	net0261#11	gnd!#1	2.592E-16
C288	net0339#2	net0346#3	2.306E-17
C289	gnd!#17	net0286#7	1.151E-16
C290	Qbar#3	net0255#6	2.041E-16
C291	net0261#10	gnd!#1	3.887E-16
C292	Q#4	net0261#9	1.396E-16
C293	net0286#6	net0187#9	1.203E-16
C294	net0346#6	gnd!#1	2.066E-17
C295	net0261#12	Qbar#3	3.155E-17
C296	net0283#4	vdd!#13	1.245E-16
C297	net0187#9	vdd!#19	3.483E-17
C298	net0286#5	net0132#5	9.049E-18
C299	net0286#6	net0132#6	5.069E-17
C300	gnd!#16	net076#4	1.159E-16
C301	phi1#8	net0255#4	1.811E-17
C302	vdd!#16	net0339#3	3.049E-16
C303	net0346#3	net076#3	1.233E-17
C304	net0283#5	net0211#6	8.709E-17
C305	net0220#7	gnd!#18	9.854E-17
C306	phi2#4	net0187#10	4.276E-17
C307	net076#6	phi1#1	1.173E-16
C308	D#1	phi2#1	4.030E-17
C309	net0286#5	net0130#9	1.134E-16
C310	gnd!#13	net0255#6	1.719E-16
C311	net0187#3	net0211#2	2.669E-16
C312	net0261#8	gnd!#1	2.621E-16
C313	vdd!#17	net0132#5	1.471E-16
C314	vdd!#4	net0261#6	7.941E-17
C315	net076#5	vdd!#2	4.526E-17
C316	net0346#3	net0130#8	2.568E-17
C317	gnd!#2	net0255#7	4.054E-17
C318	gnd!#8	net0286#7	4.249E-17
C319	net0261#5	gnd!#1	1.741E-16
C320	D#1	net0220#7	4.971E-17
C321	net0261#4	gnd!#1	7.760E-17
C322	net076#5	phi1#3	4.257E-17
C323	gnd!#3	net0261#3	3.547E-17
C324	net0130#2	net0132#6	5.148E-17
C325	net0220#5	gnd!#1	1.084E-16
C326	gnd!#6	net0130#6	5.898E-17
C327	net0339#3	net076#2	3.940E-17
C328	net0132#3	vdd!#2	2.145E-17
C329	gnd!#8	net0132#4	1.501E-16
C330	Qbar#3	gnd!#1	1.276E-16
C331	gnd!#14	net0346#7	1.151E-16
C332	net0132#5	net0130#8	1.798E-17
C333	Q#3	net0255#6	1.802E-17
C334	Q#2	net0261#10	7.559E-17
C335	net076#7	gnd!#15	1.281E-16
C336	net0346#5	net0261#6	2.351E-16
C337	gnd!#13	net0261#12	6.303E-17
C338	Qbar#3	net0261#10	7.639E-18
C339	D#2	net0220#7	1.939E-17
C340	net0187#3	net0211#6	9.562E-17
C341	net0286#6	net0220#5	2.811E-16
C342	gnd!#13	net0261#11	7.867E-17
C343	net0187#9	net0130#2	3.108E-17
C344	phi1#6	net0183#9	1.805E-17
C345	D#1	phi2#2	1.331E-17
C346	net0255#8	gnd!#1	4.653E-16
C347	net0211#2	gnd!#1	7.461E-16
C348	net0339#6	net076#5	3.667E-17
C349	gnd!#16	net076#2	4.927E-17
C350	net0286#6	phi2#4	4.362E-17
C351	gnd!#9	net0132#4	1.850E-16
C352	vdd!#10	net0187#12	8.206E-17
C353	net0255#4	gnd!#1	4.695E-16
C354	vdd!#14	net0261#6	1.473E-16
C355	net0220#5	gnd!#19	5.152E-17
C356	net0261#2	gnd!#1	7.202E-17
C357	net0339#5	net076#6	4.382E-17
C358	net0187#3	net0211#3	7.752E-17
C359	gnd!#19	D#1	2.549E-16
C360	net0130#3	net0286#7	1.391E-17
C361	vdd!#16	net076#2	8.617E-17
C362	gnd!#3	net0255#7	2.411E-16
C363	Qbar#2	net0255#6	1.175E-16
C364	vdd!#4	net0255#9	7.935E-17
C365	Q#3	net0261#11	7.762E-17
C366	net0346#5	net0255#9	1.209E-17
C367	gnd!#13	net0261#10	3.319E-17
C368	net0220#7	gnd!#1	7.930E-18
C369	net076#7	phi1#3	2.518E-17
C370	net0130#4	net0132#5	2.600E-17
C371	phi2#3	net0187#12	1.737E-17
C372	net0183#6	net076#6	2.048E-17
C373	net0183#11	gnd!#1	5.649E-16
C374	net076#2	phi1#5	7.615E-17
C375	phi1#8	net076#6	4.094E-17
C376	net0261#12	net0255#6	3.010E-17
C377	net0339#5	vdd!#2	1.144E-16
C378	phi1#3	net0183#9	4.056E-17
C379	net0261#12	Q#3	1.920E-16
C380	gnd!#6	phi1#5	3.098E-16
C381	net076#6	net0183#3	1.212E-16
C382	net0130#2	net0132#5	1.455E-16
C383	net0220#6	vdd!#18	1.598E-16
C384	net0283#2	vdd!#13	1.770E-16
C385	vdd!#14	net0255#9	1.471E-16
C386	net0187#5	net0211#2	6.701E-17
C387	Q#1	net0255#6	6.686E-18
C388	net0132#3	net0187#12	1.354E-16
C389	net0211#5	vdd!#11	1.002E-16
C390	net0339#4	vdd!#7	6.378E-17
C391	D#2	gnd!#19	4.058E-17
C392	phi2#6	net0211#3	4.968E-17
C393	net0220#5	net0187#10	1.216E-17
C394	net0183#5	net076#6	1.140E-17
C395	phi2#6	net0187#3	8.126E-17
C396	vdd!#16	net0346#2	5.016E-17
C397	vdd!#10	phi2#3	7.475E-17
C398	net0346#5	vdd!#4	8.758E-17
C399	Q#3	net0261#10	8.053E-17
C400	net0183#6	net076#7	3.846E-17
C401	phi1#4	gnd!#1	1.617E-15
C402	vdd!#17	net0130#9	3.409E-17
C403	net0339#5	net076#5	3.251E-16
C404	phi2#5	gnd!#1	1.446E-15
C405	phi1#1	gnd!#1	3.709E-17
C406	net076#5	vdd!#5	7.593E-17
C407	vdd!#2	net0130#7	2.645E-16
C408	net0132#6	net0130#9	2.525E-17
C409	net0187#6	gnd!#1	1.204E-16
C410	net0183#5	net0339#6	3.582E-17
C411	vdd!#18	net0187#12	1.224E-16
C412	net0220#5	phi2#4	1.644E-16
C413	net0346#7	net0261#8	7.831E-17
C414	net0130#4	net0286#5	9.345E-17
C415	vdd!#5	net0183#8	8.206E-17
C416	net0187#7	net0283#5	1.758E-16
C417	net0220#4	phi2#6	1.790E-17
C418	gnd!#6	net076#4	9.108E-17
C419	Q#1	net0346#5	1.583E-17
C420	net0220#5	net0211#6	1.204E-16
C421	net0132#3	phi2#3	1.082E-17
C422	phi2#7	net0211#4	1.897E-17
C423	net0130#6	gnd!#1	9.296E-16
C424	net0339#6	net0183#7	7.847E-17
C425	net0183#7	vdd!#2	1.144E-16
C426	net076#2	gnd!#1	4.364E-16
C427	net0283#6	vdd!#2	7.240E-17
C428	net0346#6	Q#3	2.941E-17
C429	net0130#3	gnd!#17	1.151E-16
C430	net0187#9	phi2#3	2.619E-17
C431	net076#6	gnd!#1	1.503E-16
C432	net0283#3	phi2#6	5.674E-18
C433	gnd!#14	net0261#8	8.103E-17
C434	vdd!#2	phi1#7	3.365E-17
C435	net0220#5	D#4	3.184E-17
C436	gnd!#9	phi2#2	1.046E-17
C437	Q#3	gnd!#1	5.631E-17
C438	net0220#3	phi2#7	1.826E-17
C439	net0286#7	net0130#10	1.367E-16
C440	net0286#4	net0220#4	2.152E-17
C441	vdd!#15	net0183#8	1.223E-16
C442	vdd!#18	phi2#3	1.480E-16
C443	net0286#2	net0220#2	8.813E-17
C444	net0220#5	phi2#3	1.186E-17
C445	net0130#2	net0286#5	1.167E-17
C446	gnd!#12	phi2#6	2.875E-16
C447	net0183#5	net0339#5	2.346E-16
C448	gnd!#19	net0220#7	2.232E-17
C449	net0346#6	net0255#8	4.452E-17
C450	net0261#3	gnd!#14	1.151E-16
C451	vdd!#11	D#5	8.342E-17
C452	phi1#5	gnd!#1	1.352E-15
C453	net0132#3	vdd!#10	7.134E-17
C454	net0211#2	D#4	7.553E-18
C455	net0346#2	gnd!#1	3.408E-16
C456	D#2	phi2#1	3.774E-17
C457	net0130#4	vdd!#17	9.211E-17
C458	net0183#3	net076#7	6.784E-17
C459	net0261#4	net0255#8	1.962E-17
C460	vdd!#5	phi1#6	8.117E-17
C461	gnd!#6	net0346#4	7.857E-17
C462	net0286#3	net0220#3	1.234E-17
C463	gnd!#14	net0255#8	7.627E-17
C464	net0220#6	phi2#3	2.623E-16
C465	net0255#4	gnd!#3	2.751E-17
C466	gnd!#17	net0130#10	9.858E-17
C467	Q#4	vdd!#2	1.187E-16
C468	gnd!#13	Qbar#3	9.850E-17
C469	net0283#6	net0211#5	3.599E-17
C470	net0261#2	net0255#8	1.802E-16
C471	net0183#5	net0339#4	7.987E-18
C472	net0346#5	net0261#7	2.057E-17
C473	net0286#7	net0346#2	9.850E-18
C474	net076#4	gnd!#1	3.677E-16
C475	vdd!#15	phi1#6	1.451E-16
C476	net0339#2	vdd!#7	6.686E-17
C477	D#2	net0220#5	1.066E-17
C478	gnd!#4	net0255#4	1.672E-16
C479	gnd!#14	net0261#5	1.322E-17
C480	net0183#6	gnd!#1	1.105E-16
C481	net0261#3	net0255#8	8.614E-17
C482	gnd!#12	net0220#4	2.059E-16
C483	Q#3	net0255#7	1.775E-17
C484	net0286#6	net0130#3	1.076E-16
C485	net076#5	phi1#6	2.243E-16
C486	net0346#7	gnd!#1	3.638E-17
C487	Qbar#2	net0255#5	1.660E-16
C488	Q#2	Qbar#2	9.872E-18
C489	net0261#4	net0346#7	9.295E-17
C490	gnd!#8	net0130#3	3.549E-17
C491	gnd!#10	D#1	1.117E-16
C492	net0339#6	vdd!#2	7.240E-17
C493	net0187#6	net0211#3	5.391E-17
C494	net0211#6	gnd!#1	5.034E-17
C495	net0346#5	Q#2	1.108E-16
C496	net0255#6	net0261#11	5.328E-17
C497	phi1#6	net0183#10	5.087E-17
C498	gnd!#17	net0132#6	1.157E-16
C499	gnd!#2	net0255#6	1.665E-16
C500	gnd!#18	phi2#5	5.943E-17
C501	net0346#4	gnd!#1	4.860E-16
C502	net0339#5	phi1#6	8.746E-18
C503	Q#1	net0255#5	2.365E-17
C504	net0187#5	D#5	3.518E-17
C505	net0132#4	gnd!#1	9.401E-16
C506	net0283#4	vdd!#2	4.930E-17
C507	phi1#1	net0183#11	2.567E-17
C508	net0283#6	net0211#4	1.623E-17
C509	net0346#7	net0261#7	5.122E-17
C510	gnd!#2	Q#3	3.547E-17
C511	phi2#4	net0187#8	2.682E-17
C512	net076	net0260	4.867E-17
C513	net0346	net076#2	5.715E-17
C514	phi2#6	net0208	2.121E-16
C515	net0286	net0187#2	1.126E-17
C516	net0286	net0211#6	1.289E-16
C517	net0187	gnd!#1	1.251E-17
C518	net0346	net0339	7.262E-17
C519	net0208	net0220#4	2.336E-18
C520	net0220#5	net0286	1.996E-16
C521	net0183#6	net0260	1.860E-16
C522	net0220	gnd!#1	5.280E-17
C523	net0339	vdd!#16	3.096E-16
C524	net0286	phi2#6	2.795E-17
C525	net0261	vdd!#4	1.191E-16
C526	Q	Qbar	1.226E-15
C527	D	phi2	1.270E-15
C528	phi2	net0132#4	7.349E-18
C529	net0187	net0286#2	3.957E-17
C530	net0183#6	net076	3.983E-17
C531	net0286	net0283#5	4.414E-17
C532	net0211	gnd!#1	6.448E-16
C533	net0183#10	net0255	5.976E-17
C534	net0286#6	net0132	1.426E-16
C535	net0286	phi2#7	2.765E-17
C536	net0187#6	net0211	1.073E-16
C537	net0286#7	net0183	9.559E-17
C538	net0268	net076#4	1.123E-16
C539	net0346	net0339#3	4.968E-17
C540	vdd!#15	net0255	1.849E-16
C541	Q	vdd!	9.784E-17
C542	net0255	net0261#2	3.563E-17
C543	net0286	net0211#2	2.669E-17
C544	net0261	net0346#5	2.725E-17
C545	net0286	net0187#3	3.424E-17
C546	gnd!#12	net0216	2.476E-16
C547	net0268	net0346#4	1.356E-16
C548	net0260	net0183#3	1.503E-16
C549	vdd!	gnd!#1	2.054E-16
C550	net0132	net0187#10	1.840E-16
C551	net0255	net0183#9	1.697E-16
C552	Qbar	vdd!	3.666E-16
C553	net0286#5	net0339	1.027E-16
C554	net0132	net0130#3	2.604E-16
C555	net0220	net0286	4.219E-16
C556	net0183#12	net0255	1.097E-16
C557	gnd!#10	net0211	9.936E-17
C558	vdd!	Qbar#1	2.685E-16
C559	net0216	net0220#4	1.123E-16
C560	net0132	net0130#2	3.484E-17
C561	net0187	gnd!#12	3.272E-16
C562	net0130	vdd!#2	1.191E-16
C563	net0255	vdd!#5	1.121E-16
C564	net0260	net0130#6	1.414E-16
C565	net0132	phi2#4	1.488E-17
C566	net076#5	net0255	1.360E-17
C567	net0216	net0286#4	1.426E-16
C568	gnd!#17	net0183	1.379E-17
C569	net0261	vdd!#14	1.849E-16
C570	net0286#6	net0346	1.008E-16
C571	Q#1	vdd!	5.120E-17
C572	phi2	gnd!#1	5.752E-17
C573	phi1#5	net0260	2.119E-16
C574	net0346	vdd!#16	4.477E-17
C575	phi1	net0255	8.231E-17
C576	net0187	net0220	1.422E-17
C577	net076	net0346#2	1.926E-17
C578	net0286	net0283	7.733E-17
C579	net0183	net076#4	1.052E-17
C580	phi1	net0261	1.147E-17
C581	vdd!	net0255#5	2.219E-16
C582	net0346	net0183#12	9.255E-18
C583	Qbar	gnd!#1	4.667E-16
C584	net0208	net0187#3	1.502E-16
C585	net0260	net076#4	2.336E-18
C586	net0187	net0220#4	1.214E-17
C587	gnd!#16	net0260	1.636E-16
C588	net0130	vdd!#17	1.849E-16
C589	net0220	net0286#2	2.155E-17
C590	net0346	net0130#6	1.066E-17
C591	net0261	net0346#6	1.000E-17
C592	net0132	net0187#8	6.029E-17
C593	net0187#6	net0208	1.828E-16
C594	net0211	gnd!#19	4.830E-17
C595	vdd!	net0261#9	1.551E-16
C596	net0286	net0187#5	2.297E-16
C597	phi2	gnd!#18	4.735E-17
C598	net0183	net0346#4	1.690E-16
C599	net0339	net0346#2	1.008E-16
C600	net0283	net0220#3	4.837E-18
C601	phi2	vdd!#18	5.981E-17
C602	gnd!#18	net0132	1.246E-16
C603	net076	net0183#3	6.457E-17
C604	net0220	net0211#2	4.761E-17
C605	Qbar	gnd!#13	3.916E-17
C606	net0286	net0283#3	5.178E-17
C607	phi2	net0220#7	7.819E-17
C608	net0283	net0286#2	1.014E-16
C609	net0346	phi1#5	2.703E-17
C610	net0187	net0286#4	1.779E-16
C611	net0220#5	net0132	1.611E-17
C612	gnd!#12	net0208	1.765E-16
C613	net0283	net0286#3	2.240E-16
C614	net0220	net0187#3	1.618E-16
C615	phi2	net0220#6	1.378E-16
C616	net0346	net076#6	2.575E-16
C617	Q#4	vdd!	1.408E-16
C618	net076	gnd!#1	7.741E-17
C619	phi2	gnd!#9	3.735E-16
C620	net0130	net0132#5	1.664E-16
C621	net0183	gnd!#1	1.686E-17
C622	net0346	net0183#2	1.161E-17
C623	net0183#12	net0261	3.234E-17
C624	net0211	D#4	1.890E-17
C625	net076	net0130#6	1.085E-17
C626	Qbar	net0261#12	2.617E-17
C627	net0132	gnd!#1	9.116E-17
C628	net0286	net0220#2	6.297E-17
C629	gnd!#6	net0260	6.865E-17
C630	Qbar	Q#1	3.087E-17
C631	net0339	net076#3	4.747E-18
C632	net0183	gnd!#16	6.990E-17
C633	net0132#3	net0130	2.272E-16
C634	net0286	vdd!#13	4.831E-17
C635	net0208	net0211#2	2.167E-17
C636	net0339	net0346#3	2.236E-16
C637	net0183	net0346	2.095E-17
C638	net076	phi1#5	5.387E-17
C639	net0283	vdd!#13	4.240E-16
C640	net0220	net0208	4.870E-17
C641	gnd!#6	net0183	1.806E-16
C642	net0286#6	net0339	3.049E-17
C643	net0346	net0130#7	1.175E-17
C644	phi2	net0286#6	1.182E-16
C645	net0339	net0130#8	6.057E-18
C646	phi2#5	net0211	1.878E-17
C647	phi2#6	net0211	1.067E-17
C648	net0183	net0346#2	4.733E-17
C649	net0220	phi2#6	5.440E-17
C650	net0183	net076	2.123E-17
C651	net0183	net0268	3.059E-16
C652	net0346	net0183#5	1.634E-16
C653	net0187#3	net0211	4.253E-17
C654	net0268	gnd!#16	1.635E-16
C655	net0346	net0339#5	4.211E-17
C656	Qbar	gnd!#2	7.224E-17
C657	net0286	net0187#9	9.772E-18
C658	net0268	net076#2	2.941E-17
C659	net0255	net0183#8	1.353E-16
C660	net0346	net0268	2.368E-17
C661	net076	gnd!#16	8.777E-17
C662	net0346	phi1#7	3.001E-17
C663	phi2	net0187#9	1.187E-16
C664	net0216	net0220#2	2.944E-17
C665	net0286	D#4	2.702E-17
C666	gnd!#6	net0268	8.405E-17
C667	phi2	vdd!#10	3.466E-16
C668	net0268	net0346#2	6.996E-18
C669	net0211	D#1	4.495E-17
C670	net076	net0268	2.238E-17
C671	net076	net0346	3.239E-16
C672	net0261	net0255#9	2.699E-16
C673	Q#2	vdd!	1.713E-17
C674	net0187#6	net0220	5.852E-17
C675	net0187	net0216	3.098E-16
C676	gnd!#8	net0183	8.019E-17
C677	phi2	net0220#5	1.341E-16
C678	Qbar	net0255#6	1.792E-17
C679	net0220	gnd!#12	8.840E-17
C680	net0346	net0183#3	3.876E-17
C681	net0339	vdd!#7	1.144E-16
C682	phi2	D#2	4.202E-17
C683	net0183	net0132#4	3.076E-17
C684	net0208	net0211#3	1.193E-16
C685	net0255	net0261	3.517E-16
C686	net0255#4	gnd!#14	9.434E-18
C687	net0261#3	gnd!#1	8.098E-18
C688	gnd!#3	net0261#8	8.425E-18
C689	net0187#7	net0220#3	3.048E-18
C690	net0220#7	net0187#10	3.514E-18
C691	net0187#5	net0220#2	4.500E-18
C692	gnd!#12	net0211#3	6.834E-18
C693	gnd!#16	net0346#4	4.595E-18
C694	net0261#3	net0183#11	4.968E-18
C695	net0261	net0183#9	7.113E-18
C696	net0261	net0183#8	7.591E-18
C697	D	net0211	4.726E-18
C698	net0211#6	D#5	6.566E-18
C699	Q#2	net0255#6	5.154E-18
C700	net0346#6	net0261#5	5.641E-18
C701	Qbar#2	net0261#9	3.591E-18
C702	net0346	net0130#9	5.710E-18
C703	net0255	phi1#3	4.998E-18
C704	net0255	phi1#6	6.171E-18
C705	net0255#2	phi1#3	9.532E-18
C706	phi1	net0255#8	9.917E-18
C707	phi1#8	net0183#10	5.847E-18
C708	phi1	net0183#7	7.766E-18
C709	net0183#5	phi1#5	7.810E-18
C710	phi2	net0132	4.077E-18
C711	phi2#5	net0132#4	4.943E-18
C712	net0130	net0187#12	7.249E-18
C713	net0130#2	net0187#8	8.422E-18
C714	net0286#7	net0132#6	6.802E-18
C715	net076#6	net0183#11	2.885E-18
C716	net0183#7	net076#3	3.048E-18
C717	net0183#5	net076#2	4.733E-18
C718	net076#6	net0183#9	5.683E-18
C719	net076#5	net0183#9	5.960E-18
C720	phi2#5	net0187#10	4.333E-18
C721	net0187#5	phi2#6	7.810E-18
C722	net0187#12	net0132#5	3.023E-18
C723	net0261#10	net0255#5	5.585E-18
C724	net0261#3	net0255#4	6.737E-18
C725	net0261#2	net0255#7	7.945E-18
C726	net0261#4	net0255#7	8.422E-18
C727	net0261#2	net0255#9	9.081E-18
C728	D	gnd!	8.601E-17
C729	Q	gnd!	4.743E-17
C730	Qbar	gnd!	2.519E-16
C731	phi1	gnd!	5.661E-17
C732	phi2	gnd!	3.250E-17
C733	net0208	gnd!	5.783E-17
C734	net0216	gnd!	4.677E-18
C735	net0268	gnd!	4.642E-18
C736	net0260	gnd!	7.676E-18
C737	net0339	gnd!	2.717E-18
C738	vdd!	gnd!	3.210E-15
C739	net0283	gnd!	2.735E-18
C740	net0255	gnd!	1.653E-16
C741	net0261	gnd!	1.419E-16
C742	net0130	gnd!	2.170E-17
C743	net0132	gnd!	9.716E-17
C744	net0211	gnd!	5.989E-19
C745	net0183	gnd!	1.498E-18
C746	net0346	gnd!	1.501E-16
C747	net076	gnd!	7.471E-18
C748	net0220	gnd!	7.675E-18
C749	net0286	gnd!	2.421E-16
C750	net0187	gnd!	5.901E-18
C751	net0255#5	gnd!	9.057E-16
C752	net0261#9	gnd!	9.435E-16
C753	net0261#6	gnd!	9.963E-16
C754	net0255#9	gnd!	1.070E-15
C755	net0183#8	gnd!	4.752E-16
C756	phi1#6	gnd!	8.070E-16
C757	net0130#7	gnd!	1.804E-15
C758	phi1#7	gnd!	8.713E-16
C759	net076#3	gnd!	6.024E-16
C760	net0346#3	gnd!	5.831E-16
C761	net0130#8	gnd!	1.490E-15
C762	net0132#5	gnd!	1.047E-15
C763	net0187#12	gnd!	4.745E-16
C764	phi2#3	gnd!	9.666E-16
C765	D#5	gnd!	1.146E-15
C766	net0211#4	gnd!	8.098E-16
C767	phi2#7	gnd!	8.825E-16
C768	net0220#3	gnd!	6.044E-16
C769	net0286#3	gnd!	5.745E-16
C770	net0255#6	gnd!	3.801E-16
C771	net0261#11	gnd!	8.274E-18
C772	net0261#8	gnd!	2.963E-18
C773	net0255#8	gnd!	4.422E-16
C774	net0183#11	gnd!	9.292E-17
C775	phi1#4	gnd!	6.361E-18
C776	net0130#6	gnd!	1.917E-16
C777	phi1#5	gnd!	2.494E-16
C778	net0346#4	gnd!	3.539E-18
C779	net0130#10	gnd!	1.110E-16
C780	net0132#6	gnd!	4.347E-16
C781	net0187#10	gnd!	7.893E-17
C782	phi2#4	gnd!	3.976E-16
C783	D#4	gnd!	5.493E-16
C784	net0211#3	gnd!	5.564E-17
C785	phi2#6	gnd!	4.012E-16
C786	net0286#4	gnd!	3.615E-18
C787	net0261#10	gnd!	5.870E-16
C788	net0261#5	gnd!	1.488E-19
C789	net0255#4	gnd!	4.522E-18
C790	net0183#10	gnd!	1.811E-16
C791	net076#2	gnd!	4.820E-16
C792	net0346#2	gnd!	8.221E-16
C793	net0130#5	gnd!	1.533E-16
C794	net0187#8	gnd!	1.099E-15
C795	phi2#2	gnd!	9.283E-20
C796	D#1	gnd!	6.700E-18
C797	net0220#2	gnd!	4.756E-16
C798	net0286#2	gnd!	7.717E-16
C799	Qbar#2	gnd!	3.156E-16
C800	net0261#12	gnd!	4.904E-18
C801	Q#1	gnd!	3.732E-17
C802	net0346#6	gnd!	3.338E-16
C803	net0261#2	gnd!	1.409E-16
C804	net0183#12	gnd!	8.783E-17
C805	phi1#1	gnd!	7.949E-18
C806	net076#6	gnd!	1.298E-16
C807	net0339#6	gnd!	3.691E-18
C808	net0183#6	gnd!	1.017E-18
C809	net0183#5	gnd!	6.354E-17
C810	net0339#4	gnd!	1.929E-18
C811	net0339#2	gnd!	8.953E-18
C812	net0286#6	gnd!	5.597E-16
C813	net0130#4	gnd!	4.184E-17
C814	net0130#2	gnd!	2.033E-16
C815	net0187#9	gnd!	1.591E-16
C816	phi2#1	gnd!	1.487E-17
C817	net0220#5	gnd!	1.002E-16
C818	D#2	gnd!	4.645E-18
C819	net0283#6	gnd!	3.691E-18
C820	net0187#6	gnd!	1.178E-16
C821	net0187#5	gnd!	1.071E-16
C822	net0283#2	gnd!	8.133E-17
C823	phi1#8	gnd!	4.548E-18
C824	Qbar#1	gnd!	6.118E-17
C825	vdd!#2	gnd!	3.165E-15
C826	Qbar#3	gnd!	6.964E-17
C827	Q#4	gnd!	1.340E-18
C828	Q#3	gnd!	1.537E-17
C829	net0346#5	gnd!	8.688E-17
C830	net0346#7	gnd!	1.050E-17
C831	vdd!#14	gnd!	2.847E-18
C832	net0261#3	gnd!	3.338E-18
C833	net0255#2	gnd!	9.834E-17
C834	vdd!#15	gnd!	6.235E-18
C835	net076#5	gnd!	1.255E-16
C836	net076#7	gnd!	4.032E-18
C837	net0339#5	gnd!	2.975E-18
C838	net0183#3	gnd!	4.661E-17
C839	net0339#3	gnd!	2.576E-18
C840	vdd!#16	gnd!	1.183E-17
C841	net0286#5	gnd!	1.526E-16
C842	vdd!#17	gnd!	5.363E-18
C843	net0130#3	gnd!	5.744E-17
C844	net0132#3	gnd!	1.823E-16
C845	vdd!#18	gnd!	6.771E-18
C846	net0220#7	gnd!	2.186E-18
C847	net0220#6	gnd!	9.041E-17
C848	vdd!#19	gnd!	6.346E-18
C849	net0211#5	gnd!	1.166E-16
C850	net0211#6	gnd!	1.893E-16
C851	net0283#5	gnd!	1.851E-18
C852	net0187#3	gnd!	3.816E-17
C853	net0283#3	gnd!	3.169E-18
C854	vdd!#13	gnd!	1.825E-15
C855	net0211#2	gnd!	3.706E-16
C856	phi2#5	gnd!	3.491E-18
C857	net0130#9	gnd!	7.743E-16
C858	phi1#3	gnd!	5.987E-16
C859	net0183#9	gnd!	8.973E-16
C860	net0261#7	gnd!	6.774E-16
C861	Q#2	gnd!	2.832E-16
C862	net0255#7	gnd!	5.379E-18
C863	vdd!#4	gnd!	1.072E-15
C864	vdd!#5	gnd!	1.068E-15
C865	vdd!#7	gnd!	1.003E-15
C866	vdd!#8	gnd!	7.927E-16
C867	vdd!#10	gnd!	1.011E-15
C868	vdd!#11	gnd!	1.106E-15
*
*
.ENDS zxw_dff
*
